-- vhdl pipelined processor