library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ALU is
port (
	A_in : in std_logic_vector (31 downto 0);
	B_in : in std_logic_vector (31 downto 0);
	opCode : in std_logic_vector (4 downto 0);
	C_out : out std_logic_vector (31 downto 0)
);
end ALU;



architecture ALU_arch of ALU is

signal hi, lo, remain_div, result_div : std_logic_vector (31 downto 0);
signal result_mult : std_logic_vector (63 downto 0);

begin

process (A_in, B_in, opCode)
begin


	case opCode is
		
		-- ADD
		when "00000" =>
			C_out <= std_logic_vector( to_unsigned( to_integer(unsigned(A_in)) + to_integer(unsigned(B_in)), C_out'length ) );


		-- SUB
		when "00001" =>
			C_out <= std_logic_vector( to_unsigned( to_integer(unsigned(A_in)) - to_integer(unsigned(B_in)), C_out'length ) );


		-- ADDI (B_in set in sign extend)
		when "00010" =>
			C_out <= std_logic_vector( to_unsigned( to_integer(unsigned(A_in)) + to_integer(unsigned(B_in)), C_out'length ) );


		-- MULT
		when "00011" =>
			result_mult <= std_logic_vector( to_unsigned( to_integer(unsigned(A_in)) * to_integer(unsigned(B_in)), 64 ) );		--32b * 32b = 64b 
			hi <= result_mult (63 downto 32);	-- 32 MSB from 64bit mult result (overflow)
			lo <= result_mult (31 downto 0);	-- 32 LSB from 64bit mult result
			C_out <= std_logic_vector( to_unsigned( to_integer(unsigned(A_in)) * to_integer(unsigned(B_in)), C_out'length ) );	-- regular multiply cast to 32 bits



		-- DIV
		when "00100" =>
			result_div <= std_logic_vector( to_unsigned( to_integer(unsigned(A_in)) / to_integer(unsigned(B_in)), C_out'length ) );		-- division result
			remain_div <= std_logic_vector( to_unsigned( to_integer(unsigned(A_in)) mod to_integer(unsigned(B_in)), remain_div'length ) );	-- remainder of division
			hi <= remain_div;		-- from MIPS reference
			lo <= result_div;		-- from MIPS reference
			C_out <= result_div;		-- output = result 



		-- SLT (set less than)
		when "00101" =>
			if (unsigned(A_in) < unsigned(B_in)) then
				C_out <= x"00000001";	-- True
			else
				C_out <= x"00000000";	-- False
			end if;


		-- SLTI (set less than immediate)  (B_in set in sign extend)
		when "00110" =>
			if (unsigned(A_in) < unsigned(B_in)) then
				C_out <= x"00000001";	-- True
			else
				C_out <= x"00000000";	-- False
			end if;



		-- AND
		when "00111" => 
			C_out <= A_in and B_in;



		-- OR
		when "01000" => 
			C_out <= A_in or B_in;


		-- NOR
		when "01001" => 
			C_out <= A_in nor B_in;


		-- XOR
		when "01010" => 
			C_out <= A_in xor B_in;


		-- ANDI  (B_in set in sign extend)
		when "01011" => 
			C_out <= A_in and B_in;


		-- ORI  (B_in set in sign extend)
		when "01100" => 
			C_out <= A_in or B_in;


		-- XORI  (B_in set in sign extend)
		when "01101" => 
			C_out <= A_in xor B_in;


		-- MFHI (move from hi)
		when "01110" => 
			C_out <= hi;	-- output saved result from MSB of mult or remainder of div


		-- MFLO (move from lo)
		when "01111" => 
			C_out <= lo;	-- output saved result from LSB of mult or result of div


		-- LUI (load upper immediate)
		when "10000" => 
			C_out <= B_in(15 downto 0) & std_logic_vector(to_unsigned(0,16));	-- output mask x11110000 (keep only 16 MSB)


		-- SLL (shift left logical)
		when "10001" =>
			C_out <= A_in((31 - to_integer(unsigned(B_in(10 downto 6)))) downto 0)  &  std_logic_vector(to_unsigned(0, to_integer(unsigned(B_in(10 downto 6)))));
			-- Shifts A left by shamt(found in B at bits 10 downto 6) 



		-- SRL (shift right logical)
		when "10010" =>
			C_out <= std_logic_vector(to_unsigned(0, to_integer(unsigned(B_in(10 downto 6)))))  &   A_in(31 downto (0 + to_integer(unsigned(B_in(10 downto 6)))));
			-- Shifts A right by shamt(found in B at bits 10 downto 6) 



		-- SRA (shift right arithmetic)
		when "10011" =>
			if A_in(31) = '0' then
				C_out <= std_logic_vector(to_unsigned(0, to_integer(unsigned(B_in(10 downto 6)))))  &   A_in(31 downto (0 + to_integer(unsigned(B_in(10 downto 6)))));
				-- add 0s at beginning (positive num)
			else
				C_out <= std_logic_vector(to_unsigned(1, to_integer(unsigned(B_in(10 downto 6)))))  &   A_in(31 downto (0 + to_integer(unsigned(B_in(10 downto 6)))));
				-- add 1s at beginning (negative num)
			end if;



		-- LW (load word)  (B_in set in sign extend)
		when "10100" =>
			C_out <= std_logic_vector( to_unsigned( to_integer(unsigned(A_in)) + to_integer(unsigned(B_in)), C_out'length ) );


		-- SW (store word)  (B_in set in sign extend)
		when "10101" =>
			C_out <= std_logic_vector( to_unsigned( to_integer(unsigned(A_in)) + to_integer(unsigned(B_in)), C_out'length ) );


		-- BEQ (branch if equal)  (condition checked in "zero?")
		when "10110" =>
			C_out <= std_logic_vector( to_unsigned(  (to_integer(unsigned(A_in)) + to_integer(unsigned(B_in)) * 4), C_out'length ) );


		-- BNE (branch if not equal)  (condition checked in "zero?")
		when "10111" =>
			C_out <= std_logic_vector( to_unsigned(  (to_integer(unsigned(A_in)) + to_integer(unsigned(B_in)) * 4), C_out'length ) );


		-- J (assume that B_in is 26 bits, LSB)
		when "11000" =>
			C_out <= A_in(31 downto 28) & B_in(25 downto 0) & "00";


		-- JR (jump register)
		when "11001" =>
			C_out <= A_in;


		-- JAL (jump and link)
		when "11010" =>
			C_out <= A_in(31 downto 28) & B_in(25 downto 0) & "00";


		when others =>
			null;

	end case;
end process;

end ALU_arch;


