-- ALU Operations